-- VHDL file
--
-- Autor: Jassan, Joel
-- Date: (mmm/YYYY)
-- 
-- Proyect Explanation:
--
--
-- Copyright 2023, Joel Jassan <joeljassan@hotmail.com>
-- All rights reserved.
---------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity ent is
	
	generic (

    );

	port (
        --input ports
		clk		  	: in std_logic;
		reset	  	: in std_logic;
		enable		: in std_logic;

        --output ports
    
    );

end entity;

architecture a_ent of ent is

    ----- Typedefs --------------------------------------------------------------------------------
    
    ----- Constants -------------------------------------------------------------------------------

    ----- Signals (i: entrada, o:salida, s:señal intermedia)---------------------------------------


begin
    ----- Components ------------------------------------------------------------------------------

    ----- Codigo ----------------------------------------------------------------------------------
    
    -- Logica Estado Siguiente

    -- Logica Salida

    
end architecture ; 
